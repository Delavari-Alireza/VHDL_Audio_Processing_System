LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;

ENTITY PROZHE IS
	PORT
	(	
		BCLK	: IN 	STD_LOGIC;
		Reset	: IN 	STD_LOGIC;
		
		DR		: IN 	STD_LOGIC;

		InST1	: IN 	STD_LOGIC_VECTOR(4 DOWNTO 0);
		InST2	: IN 	STD_LOGIC_VECTOR(4 DOWNTO 0);

		OutST	: IN 	STD_LOGIC_VECTOR(4 DOWNTO 0);

		DX		: OUT 	STD_LOGIC
		
	);
END PROZHE;

ARCHITECTURE behavioral OF PROZHE IS

	TYPE prom_memory_AtoL IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

	TYPE prom_memory_U2law IS ARRAY (0 TO 8191) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

	CONSTANT prom_AtoL : prom_memory_AtoL := ( "1110101010000000" , "1110101110000000" , "1110100010000000" , "1110100110000000" , "1110111010000000" , "1110111110000000" , "1110110010000000" , "1110110110000000" , "1110001010000000" , "1110001110000000" , "1110000010000000" , "1110000110000000" , "1110011010000000" , "1110011110000000" , "1110010010000000" , "1110010110000000" , "1111010101000000" , "1111010111000000" , "1111010001000000" , "1111010011000000" , "1111011101000000" , "1111011111000000" , "1111011001000000" , "1111011011000000" , "1111000101000000" , "1111000111000000" , "1111000001000000" , "1111000011000000" , "1111001101000000" , "1111001111000000" , "1111001001000000" , "1111001011000000" , "1010101000000000" , "1010111000000000" , "1010001000000000" , "1010011000000000" , "1011101000000000" , "1011111000000000" , "1011001000000000" , "1011011000000000" , "1000101000000000" , "1000111000000000" , "1000001000000000" , "1000011000000000" , "1001101000000000" , "1001111000000000" , "1001001000000000" , "1001011000000000" , "1101010100000000" , "1101011100000000" , "1101000100000000" , "1101001100000000" , "1101110100000000" , "1101111100000000" , "1101100100000000" , "1101101100000000" , "1100010100000000" , "1100011100000000" , "1100000100000000" , "1100001100000000" , "1100110100000000" , "1100111100000000" , "1100100100000000" , "1100101100000000" , "1111111010101000" , "1111111010111000" , "1111111010001000" , "1111111010011000" , "1111111011101000" , "1111111011111000" , "1111111011001000" , "1111111011011000" , "1111111000101000" , "1111111000111000" , "1111111000001000" , "1111111000011000" , "1111111001101000" , "1111111001111000" , "1111111001001000" , "1111111001011000" , "1111111110101000" , "1111111110111000" , "1111111110001000" , "1111111110011000" , "1111111111101000" , "1111111111111000" , "1111111111001000" , "1111111111011000" , "1111111100101000" , "1111111100111000" , "1111111100001000" , "1111111100011000" , "1111111101101000" , "1111111101111000" , "1111111101001000" , "1111111101011000" , "1111101010100000" , "1111101011100000" , "1111101000100000" , "1111101001100000" , "1111101110100000" , "1111101111100000" , "1111101100100000" , "1111101101100000" , "1111100010100000" , "1111100011100000" , "1111100000100000" , "1111100001100000" , "1111100110100000" , "1111100111100000" , "1111100100100000" , "1111100101100000" , "1111110101010000" , "1111110101110000" , "1111110100010000" , "1111110100110000" , "1111110111010000" , "1111110111110000" , "1111110110010000" , "1111110110110000" , "1111110001010000" , "1111110001110000" , "1111110000010000" , "1111110000110000" , "1111110011010000" , "1111110011110000" , "1111110010010000" , "1111110010110000" , "0001010110000000" , "0001010010000000" , "0001011110000000" , "0001011010000000" , "0001000110000000" , "0001000010000000" , "0001001110000000" , "0001001010000000" , "0001110110000000" , "0001110010000000" , "0001111110000000" , "0001111010000000" , "0001100110000000" , "0001100010000000" , "0001101110000000" , "0001101010000000" , "0000101011000000" , "0000101001000000" , "0000101111000000" , "0000101101000000" , "0000100011000000" , "0000100001000000" , "0000100111000000" , "0000100101000000" , "0000111011000000" , "0000111001000000" , "0000111111000000" , "0000111101000000" , "0000110011000000" , "0000110001000000" , "0000110111000000" , "0000110101000000" , "0101011000000000" , "0101001000000000" , "0101111000000000" , "0101101000000000" , "0100011000000000" , "0100001000000000" , "0100111000000000" , "0100101000000000" , "0111011000000000" , "0111001000000000" , "0111111000000000" , "0111101000000000" , "0110011000000000" , "0110001000000000" , "0110111000000000" , "0110101000000000" , "0010101100000000" , "0010100100000000" , "0010111100000000" , "0010110100000000" , "0010001100000000" , "0010000100000000" , "0010011100000000" , "0010010100000000" , "0011101100000000" , "0011100100000000" , "0011111100000000" , "0011110100000000" , "0011001100000000" , "0011000100000000" , "0011011100000000" , "0011010100000000" , "0000000101011000" , "0000000101001000" , "0000000101111000" , "0000000101101000" , "0000000100011000" , "0000000100001000" , "0000000100111000" , "0000000100101000" , "0000000111011000" , "0000000111001000" , "0000000111111000" , "0000000111101000" , "0000000110011000" , "0000000110001000" , "0000000110111000" , "0000000110101000" , "0000000001011000" , "0000000001001000" , "0000000001111000" , "0000000001101000" , "0000000000011000" , "0000000000001000" , "0000000000111000" , "0000000000101000" , "0000000011011000" , "0000000011001000" , "0000000011111000" , "0000000011101000" , "0000000010011000" , "0000000010001000" , "0000000010111000" , "0000000010101000" , "0000010101100000" , "0000010100100000" , "0000010111100000" , "0000010110100000" , "0000010001100000" , "0000010000100000" , "0000010011100000" , "0000010010100000" , "0000011101100000" , "0000011100100000" , "0000011111100000" , "0000011110100000" , "0000011001100000" , "0000011000100000" , "0000011011100000" , "0000011010100000" , "0000001010110000" , "0000001010010000" , "0000001011110000" , "0000001011010000" , "0000001000110000" , "0000001000010000" , "0000001001110000" , "0000001001010000" , "0000001110110000" , "0000001110010000" , "0000001111110000" , "0000001111010000" , "0000001100110000" , "0000001100010000" , "0000001101110000" , "0000001101010000" );

	CONSTANT prom_U2law : prom_memory_U2law := ( "11111111" , "11111110" , "11111101" , "11111100" , "11111011" , "11111010" , "11111001" , "11111000" , "11110111" , "11110110" , "11110101" , "11110100" , "11110011" , "11110010" , "11110001" , "11110000" , "11101111" , "11101111" , "11101110" , "11101110" , "11101101" , "11101101" , "11101100" , "11101100" , "11101011" , "11101011" , "11101010" , "11101010" , "11101001" , "11101001" , "11101000" , "11101000" , "11100111" , "11100111" , "11100110" , "11100110" , "11100101" , "11100101" , "11100100" , "11100100" , "11100011" , "11100011" , "11100010" , "11100010" , "11100001" , "11100001" , "11100000" , "11100000" , "11011111" , "11011111" , "11011111" , "11011111" , "11011110" , "11011110" , "11011110" , "11011110" , "11011101" , "11011101" , "11011101" , "11011101" , "11011100" , "11011100" , "11011100" , "11011100" , "11011011" , "11011011" , "11011011" , "11011011" , "11011010" , "11011010" , "11011010" , "11011010" , "11011001" , "11011001" , "11011001" , "11011001" , "11011000" , "11011000" , "11011000" , "11011000" , "11010111" , "11010111" , "11010111" , "11010111" , "11010110" , "11010110" , "11010110" , "11010110" , "11010101" , "11010101" , "11010101" , "11010101" , "11010100" , "11010100" , "11010100" , "11010100" , "11010011" , "11010011" , "11010011" , "11010011" , "11010010" , "11010010" , "11010010" , "11010010" , "11010001" , "11010001" , "11010001" , "11010001" , "11010000" , "11010000" , "11010000" , "11010000" , "11001111" , "11001111" , "11001111" , "11001111" , "11001111" , "11001111" , "11001111" , "11001111" , "11001110" , "11001110" , "11001110" , "11001110" , "11001110" , "11001110" , "11001110" , "11001110" , "11001101" , "11001101" , "11001101" , "11001101" , "11001101" , "11001101" , "11001101" , "11001101" , "11001100" , "11001100" , "11001100" , "11001100" , "11001100" , "11001100" , "11001100" , "11001100" , "11001011" , "11001011" , "11001011" , "11001011" , "11001011" , "11001011" , "11001011" , "11001011" , "11001010" , "11001010" , "11001010" , "11001010" , "11001010" , "11001010" , "11001010" , "11001010" , "11001001" , "11001001" , "11001001" , "11001001" , "11001001" , "11001001" , "11001001" , "11001001" , "11001000" , "11001000" , "11001000" , "11001000" , "11001000" , "11001000" , "11001000" , "11001000" , "11000111" , "11000111" , "11000111" , "11000111" , "11000111" , "11000111" , "11000111" , "11000111" , "11000110" , "11000110" , "11000110" , "11000110" , "11000110" , "11000110" , "11000110" , "11000110" , "11000101" , "11000101" , "11000101" , "11000101" , "11000101" , "11000101" , "11000101" , "11000101" , "11000100" , "11000100" , "11000100" , "11000100" , "11000100" , "11000100" , "11000100" , "11000100" , "11000011" , "11000011" , "11000011" , "11000011" , "11000011" , "11000011" , "11000011" , "11000011" , "11000010" , "11000010" , "11000010" , "11000010" , "11000010" , "11000010" , "11000010" , "11000010" , "11000001" , "11000001" , "11000001" , "11000001" , "11000001" , "11000001" , "11000001" , "11000001" , "11000000" , "11000000" , "11000000" , "11000000" , "11000000" , "11000000" , "11000000" , "11000000" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111111" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111110" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111101" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111100" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111011" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111010" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111001" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10111000" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110111" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110110" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110101" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110100" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110011" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110010" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110001" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10110000" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101111" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101110" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101101" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101100" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101011" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101010" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101001" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10101000" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100111" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100110" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100101" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100100" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100011" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100010" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100001" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10100000" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011111" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011110" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011101" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011100" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011011" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011010" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011001" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10011000" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010111" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010110" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010101" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010100" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010011" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010010" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010001" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10010000" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001111" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001110" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001101" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001100" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001011" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001010" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001001" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10001000" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000111" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000110" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000101" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000100" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000011" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000010" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000001" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "10000000" , "01111111" , "01110000" , "01110001" , "01110010" , "01110011" , "01110100" , "01110101" , "01110110" , "01110111" , "01111000" , "01111001" , "01111010" , "01111011" , "01111100" , "01111101" , "01111110" , "01111111" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000001" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000010" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000011" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000100" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000101" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000110" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00000111" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001000" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001001" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001010" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001011" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001100" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001101" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001110" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00001111" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010000" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010001" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010010" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010011" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010100" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010101" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010110" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00010111" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011000" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011001" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011010" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011011" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011100" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011101" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011110" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00011111" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100000" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100001" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100010" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100011" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100100" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100101" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100110" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00100111" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101000" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101001" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101010" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101011" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101100" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101101" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101110" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00101111" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110000" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110001" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110010" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110011" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110100" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110101" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110110" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00110111" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111000" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111001" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111010" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111011" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111100" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111101" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111110" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "00111111" , "01000000" , "01000000" , "01000000" , "01000000" , "01000000" , "01000000" , "01000000" , "01000000" , "01000001" , "01000001" , "01000001" , "01000001" , "01000001" , "01000001" , "01000001" , "01000001" , "01000010" , "01000010" , "01000010" , "01000010" , "01000010" , "01000010" , "01000010" , "01000010" , "01000011" , "01000011" , "01000011" , "01000011" , "01000011" , "01000011" , "01000011" , "01000011" , "01000100" , "01000100" , "01000100" , "01000100" , "01000100" , "01000100" , "01000100" , "01000100" , "01000101" , "01000101" , "01000101" , "01000101" , "01000101" , "01000101" , "01000101" , "01000101" , "01000110" , "01000110" , "01000110" , "01000110" , "01000110" , "01000110" , "01000110" , "01000110" , "01000111" , "01000111" , "01000111" , "01000111" , "01000111" , "01000111" , "01000111" , "01000111" , "01001000" , "01001000" , "01001000" , "01001000" , "01001000" , "01001000" , "01001000" , "01001000" , "01001001" , "01001001" , "01001001" , "01001001" , "01001001" , "01001001" , "01001001" , "01001001" , "01001010" , "01001010" , "01001010" , "01001010" , "01001010" , "01001010" , "01001010" , "01001010" , "01001011" , "01001011" , "01001011" , "01001011" , "01001011" , "01001011" , "01001011" , "01001011" , "01001100" , "01001100" , "01001100" , "01001100" , "01001100" , "01001100" , "01001100" , "01001100" , "01001101" , "01001101" , "01001101" , "01001101" , "01001101" , "01001101" , "01001101" , "01001101" , "01001110" , "01001110" , "01001110" , "01001110" , "01001110" , "01001110" , "01001110" , "01001110" , "01001111" , "01001111" , "01001111" , "01001111" , "01001111" , "01001111" , "01001111" , "01001111" , "01010000" , "01010000" , "01010000" , "01010000" , "01010001" , "01010001" , "01010001" , "01010001" , "01010010" , "01010010" , "01010010" , "01010010" , "01010011" , "01010011" , "01010011" , "01010011" , "01010100" , "01010100" , "01010100" , "01010100" , "01010101" , "01010101" , "01010101" , "01010101" , "01010110" , "01010110" , "01010110" , "01010110" , "01010111" , "01010111" , "01010111" , "01010111" , "01011000" , "01011000" , "01011000" , "01011000" , "01011001" , "01011001" , "01011001" , "01011001" , "01011010" , "01011010" , "01011010" , "01011010" , "01011011" , "01011011" , "01011011" , "01011011" , "01011100" , "01011100" , "01011100" , "01011100" , "01011101" , "01011101" , "01011101" , "01011101" , "01011110" , "01011110" , "01011110" , "01011110" , "01011111" , "01011111" , "01011111" , "01011111" , "01100000" , "01100000" , "01100001" , "01100001" , "01100010" , "01100010" , "01100011" , "01100011" , "01100100" , "01100100" , "01100101" , "01100101" , "01100110" , "01100110" , "01100111" , "01100111" , "01101000" , "01101000" , "01101001" , "01101001" , "01101010" , "01101010" , "01101011" , "01101011" , "01101100" , "01101100" , "01101101" , "01101101" , "01101110" , "01101110" , "01101111" , "01101111" , "01110000" , "01110001" , "01110010" , "01110011" , "01110100" , "01110101" , "01110110" , "01110111" , "01111000" , "01111001" , "01111010" , "01111011" , "01111100" , "01111101" , "01111110" );
	
	
	
	signal FS1					: STD_LOGIC;
	signal ready				: STD_LOGIC := '0';

	signal sumReady				: STD_LOGIC := '0'; 

	signal flag_EndRead1		: boolean := false;
	signal flag_EndRead2		: boolean := false;

	signal first_Wave			: STD_LOGIC_VECTOR(7 DOWNTO 0);
	signal second_Wave			: STD_LOGIC_VECTOR(7 DOWNTO 0);

	signal first_Wave_linear	: STD_LOGIC_VECTOR(15 DOWNTO 0);
	signal second_Wave_linear	: STD_LOGIC_VECTOR(15 DOWNTO 0);

	signal first_Wave_linear_int		: integer:= 0;
	signal second_Wave_linear_int		: integer:= 0;

	signal sum_Wave_int			: integer:= 0;
	signal sum_Wave				: STD_LOGIC_VECTOR(15 DOWNTO 0);

	signal out_wave				: STD_LOGIC_VECTOR(7 DOWNTO 0);

	signal clock_counter 		: integer:= 0;
	signal Courrent_TimeSlot 	: integer:= 0;

	signal InST1_integer		: integer:= 0;
	signal InST2_integer		: integer:= 0;
	signal OutST_integer		: integer:= 0;

	signal clk_1				: boolean := true;
	signal clk_2				: boolean := false;
	signal clk_3				: boolean := false;
	signal clk_4				: boolean := false;
	signal clk_5				: boolean := false;
	
	
	

BEGIN


	InST1_integer 	<= to_integer(unsigned(InST1));
	InST2_integer 	<= to_integer(unsigned(InST2));
	OutST_integer 	<= to_integer(unsigned(OutST));


	PROCESS(BCLK)
	BEGIN
		IF (BCLK = '1' AND BCLK'EVENT) THEN  -- Positive Edge
			
		    FS1 <= '0';
			clock_counter <= clock_counter + 1;

			

			Courrent_TimeSlot <= (clock_counter + 1) / 8 ;

			if (clock_counter = 255) then
				Courrent_TimeSlot <= 31;
				FS1 <= '1'; 
			elsif (clock_counter > 255) then 
				Courrent_TimeSlot <= -1;
			end if;



			

			IF (Reset = '1' ) THEN

				clock_counter <= 0;
				first_Wave <= "UUUUUUUU";
				second_Wave <= "UUUUUUUU";
				sum_Wave <= "UUUUUUUUUUUUUUUU";
				out_wave <= "UUUUUUUU";
				Courrent_TimeSlot <= 0;
				flag_EndRead1 <= false;
				flag_EndRead2 <= false;
				ready <= '0';

			END IF;

			IF ( FS1 = '1') THEN

				clock_counter <= 0;
				Courrent_TimeSlot <= 0;

			END IF;




			IF (Courrent_TimeSlot = InST1_integer) THEN

				first_Wave <= DR & first_Wave(7 downto 1) ;

				IF (clock_counter mod 8 = 7) then
					flag_EndRead1 <= true;
				end IF;	

			elsif (Courrent_TimeSlot = InST2_integer) then 

				second_Wave <= DR & second_Wave(7 downto 1);

				IF (clock_counter mod 8 = 7) then
					flag_EndRead2 <= true;
				end IF;	

			elsif (Courrent_TimeSlot = OutST_integer AND ready = '1') then 	

				DX <= out_wave(0);

				out_wave <= '0' & out_wave(7 downto 1);
				
				
				IF (clock_counter mod 8 = 7) then
					ready <= '0';

				end IF;	

			else 
				DX	<= 'Z';
			END IF;

			IF (flag_EndRead1 AND flag_EndRead2 ) THEN

				
				IF ( clk_1) THEN	--------------- To linear form --------------------
					first_Wave_linear <= prom_AtoL(CONV_INTEGER(first_Wave));

					second_Wave_linear <= prom_AtoL(CONV_INTEGER(second_Wave));

					clk_1 <= false;
					clk_2 <= true;

				elsif (clk_2) THEN	------   integer form ------

					first_Wave_linear_int 	<= to_integer(unsigned(first_Wave_linear));
					second_Wave_linear_int	<= to_integer(unsigned(second_Wave_linear));

					clk_2 <= false;
					clk_3 <= true;
				elsif (clk_3) THEN	--- SUM
					sum_Wave_int <= first_Wave_linear_int + second_Wave_linear_int;
					clk_3 <= false;
					clk_4 <= true;

				elsif (clk_4) THEN	--- SUM to vector
					sum_Wave <= std_logic_vector(to_unsigned(sum_Wave_int, sum_Wave'length));
					
					
					clk_4 <= false;
					clk_5 <= true;

				elsif (clk_5) THEN

					
					if (CONV_INTEGER(sum_wave) > 8191) then  -- NOT OK
							
						out_wave <= prom_U2law(8191); -- be khater kochaki size dade vorodi jadval

					else -- OK
						out_wave <= prom_U2law(CONV_INTEGER(sum_wave));
					end if;
					
					ready <= '1';
					flag_EndRead1 <= false;		-- baraye in ke dobar ein if ejra nashe
					flag_EndRead2 <= false;
					clk_5 <= false;
					clk_1 <= true;


			
					
				END IF;	

			END IF;
			
		END IF;
	END PROCESS;



END behavioral;